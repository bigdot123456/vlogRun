QuestaSim-64 vlog 2020.3 Compiler 2020.07 Jul 12 2020
Start time: 11:12:27 on Aug 30,2021
vlog oran_radio_if_sspuc_ti_src_hdl_noenc.sv 
-- Compiling module sspuc_ti_sv
-- Compiling module sspuc_ul_src
-- Compiling module sspuc_ul_src_bf_buf_model
** Warning: oran_radio_if_sspuc_ti_src_hdl_noenc.sv(722): (vlog-13314) Defaulting port 'cc_ul_ud_iq_width' kind to 'var' rather than 'wire' due to default compile option setting of -svinputport=relaxed.
** Warning: oran_radio_if_sspuc_ti_src_hdl_noenc.sv(723): (vlog-13314) Defaulting port 'cc_ul_ud_comp_meth' kind to 'var' rather than 'wire' due to default compile option setting of -svinputport=relaxed.
-- Compiling module sspuc_push_pull_buf
-- Compiling module sspuc_ul_prach_gen
-- Compiling module sspuc_dl_sink

Top level modules:
	sspuc_ti_sv
End time: 11:12:27 on Aug 30,2021, Elapsed time: 0:00:00
Errors: 0, Warnings: 2
