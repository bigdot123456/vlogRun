QuestaSim-64 vlog 2020.3 Compiler 2020.07 Jul 12 2020
Start time: 11:12:27 on Aug 30,2021
vlog sspuc_ti_v2sv.sv 
-- Compiling module sspuc_ti_v2sv

Top level modules:
	sspuc_ti_v2sv
End time: 11:12:27 on Aug 30,2021, Elapsed time: 0:00:00
Errors: 0, Warnings: 0
